`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////
// Module : URMTriggerTest
// Purpose: Test bench for the URMTrigger
//////////////////////////////////////////////////////////////////////////////
module URMTriggerTest;
  
//////////////////////////////////////////////////////////////////////////////
// Registers
//////////////////////////////////////////////////////////////////////////////
reg Clock;
reg TriggerIn;
 
//////////////////////////////////////////////////////////////////////////////
// Wires
//////////////////////////////////////////////////////////////////////////////
wire TriggerOut;

// Instantiate the Unit Under Test (UUT)
// Test the ultrasonic range module trigger in Verilog
URMTrigger uut
(
  .Clock(Clock), 
  .TriggerIn(TriggerIn),
  .TriggerOut(TriggerOut)
);
 
initial begin
  // Initialize Inputs
  Clock = 0;
  TriggerIn = 0;
end
 
always begin
  // Toggle the state of the clock every 10ns
  #10 Clock = !Clock;
end

always begin
  #10;
  TriggerIn = 1;
  #20;
  TriggerIn = 0;
  #100000;
end
      
endmodule


