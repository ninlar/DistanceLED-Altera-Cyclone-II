`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////
// Module : ClockDividerTest
// Purpose: Test bench for the ClockDivider
//////////////////////////////////////////////////////////////////////////////
module ClockDividerTest;
  
//////////////////////////////////////////////////////////////////////////////
// Registers
//////////////////////////////////////////////////////////////////////////////
reg ClockIn;
 
//////////////////////////////////////////////////////////////////////////////
// Wires
//////////////////////////////////////////////////////////////////////////////
wire ClockOut;

// Instantiate the Unit Under Test (UUT)
// Test the clock divider in Verilog
ClockDivider uut
(
   .ClockIn(ClockIn), 
   .ClockOut(ClockOut)
);

// Divide the clock by 50 for 1MHz
defparam uut.DIVISOR = 50;
 
initial begin
  // Initialize Inputs
  ClockIn = 0;
end
 
always begin
  // Toggle the state of the clock every 10ns
  #10 ClockIn = !ClockIn;
end
      
endmodule
